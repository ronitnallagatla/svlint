module identifier_matches_filename;
endmodule