module identifier_matches_filename;
endfunction